library verilog;
use verilog.vl_types.all;
entity procesador_tb is
end procesador_tb;
